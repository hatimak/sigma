`timescale 1ps / 1ps

module matrix_add_tb ();

    reg [255:0]  mat1_a, mat1_b;
    wire [255:0] mat1_sum;
    reg [575:0]  mat2_a, mat2_b;
    wire [575:0] mat2_sum;
    reg          rst, clk, enable1, enable2;
    wire         ready1, ready2;

    matrix_add #(.SIZE(2)) UUT_1(
        .sum    (mat1_sum),
        .ready  (ready1),
        .op_a   (mat1_a),
        .op_b   (mat1_b),
        .enable (enable1),
        .clk    (clk),
        .rst    (rst)
        );

    matrix_add #(.SIZE(3)) UUT_2(
        .sum    (mat2_sum),
        .ready  (ready2),
        .op_a   (mat2_a),
        .op_b   (mat2_b),
        .enable (enable2),
        .clk    (clk),
        .rst    (rst)
        );

    initial begin
        $dumpfile("matrix_add.vcd");
        $dumpvars(0, matrix_add_tb);
        rst = 1'b1;
        clk = 1'b0;
        enable1 = 1'b0;
        enable2 = 1'b0;
        #20000;
        rst = 1'b0;
        /* +-                                      -+   +-                                      -+   +-                                               -+
         * |  3.4500000000e+002  -9.0300000000e+002 |   | -3.4400000000e+002   2.1000000000e+001 |   | 3.422700000000000e+001  -8.820000000000000e+002 |
         * |                                        | + |                                        | = |                                                 |
         * | -1.0000000000e-309  -4.0600000000e+001 |   |  1.1000000000e-309  -3.5700000000e+001 |   | 9.999999999999969e-311  -7.630000000000001e+001 |
         * +-                                      -+   +-                                      -+   +-                                               -+
         */
        mat1_a = 256'b1100000001000100010011001100110011001100110011001100110011001101_1000000000000000101110000001010101110010011010001111110110101110_1100000010001100001110000000000000000000000000000000000000000000_0100000001110101100100000000000000000000000000000000000000000000;
        mat1_b = 256'b1100000001000001110110011001100110011001100110011001100110011010_0000000000000000110010100111110111111101110110011110001111011001_0100000000110101000000000000000000000000000000000000000000000000_1100000001110101100000000000000000000000000000000000000000000000;
        #10;
        enable1 = 1'b1;
        #5000;
        enable1 = 1'b0;
        #300000;
        $display("[a]_{2x2} + [b]_{2x2} = [c]_{2x2}");
        if (mat1_sum[63:0] == 64'h3FF0000000000000) begin
            $display($time,"ps: Pass! a_11 + b_11 = c_11 (%h)", mat1_sum[63:0]);
        end else begin
            $display($time,"ps: Error! a_11 + b_11 != c_11 (%h)", mat1_sum[63:0]);
        end
        if (mat1_sum[127:64] == 64'hC08B900000000000) begin
            $display($time,"ps: Pass! a_12 + b_12 = c_12 (%h)", mat1_sum[127:64]);
        end else begin
            $display($time,"ps: Error! a_12 + b_12 != c_12 (%h)", mat1_sum[127:64]);
        end
        if (mat1_sum[191:128] == 64'h000012688B70E62B) begin
            $display($time,"ps: Pass! a_21 + b_21 = c_21 (%h)", mat1_sum[191:128]);
        end else begin
            $display($time,"ps: Error! a_21 + b_21 != c_21 (%h)", mat1_sum[191:128]);
        end
        if (mat1_sum[255:192] == 64'hC053133333333334) begin
            $display($time,"ps: Pass! a_22 + b_22 = c_22 (%h)", mat1_sum[255:192]);
        end else begin
            $display($time,"ps: Error! a_22 + b_22 != c_22 (%h)", mat1_sum[255:192]);
        end

        /* +-                                                          -+   +-                                                          -+   +-                                                                         -+
         * |  3.0000000000e-310   4.4000000000e+001   3.9800000000e+000 |   |  4.0000000000e-304   7.9000000000e-002   3.7700000000e+000 |   |  4.000003000000000e-304   4.407900000000000e+001   7.750000000000000e+000 |
         * |  5.0000000000e-308   2.1000000000e-308   5.4000000000e+001 | + |  2.0000000000e-312   2.0000000000e-308   0.0000000000e+000 | = |  5.000199999999999e-308   4.100000000000000e-308   5.400000000000000e+001 |
         * | -4.0600000000e+001  -1.0000000000e-309   2.0000000000e-311 |   | -3.5700000000e+001   1.1000000000e-309   0.0000000000e+000 |   | -7.630000000000001e+001   9.999999999999969e-311   1.999999999999895e-311 |
         * +-                                                          -+   +-                                                          -+   +-                                                                         -+
         */
        mat2_a = 576'b0000000000000000000000111010111010000010010010011100011110100010_1000000000000000101110000001010101110010011010001111110110101110_1100000001000100010011001100110011001100110011001100110011001101_0100000001001011000000000000000000000000000000000000000000000000_0000000000001111000110011100001001100010100111001100111101010011_0000000000100001111110100001100000101100010000001100011000001101_0100000000001111110101110000101000111101011100001010001111010111_0100000001000110000000000000000000000000000000000000000000000000_0000000000000000001101110011100110100010010100101011001010000001;
        mat2_b = 576'b0000000000000000000000000000000000000000000000000000000000000000_0000000000000000110010100111110111111101110110011110001111011001_1100000001000001110110011001100110011001100110011001100110011010_0000000000000000000000000000000000000000000000000000000000000000_0000000000001110011000011010110011110000001100111101000110100100_0000000000000000000000000101111001000000001110101001001111110110_0100000000001110001010001111010111000010100011110101110000101001_0011111110110100001110010101100000010000011000100100110111010011_0000000011110001100011100011101110011011001101110100000101101001;
        #10;
        enable2 = 1'b1;
        #10000;
        enable2 = 1'b0;
        #300000;
        $display("");
        $display("[e]_{3x3} + [f]_{3x3} = [g]_{3x3}");
        if (mat2_sum[63:0] == 64'h00F18E3C781DCAB4) begin
            $display($time,"ps: Pass! e_11 + f_11 = g_11 (%h)", mat2_sum[63:0]);
        end else begin
            $display($time,"ps: Error! e_11 + f_11 != g_11 (%h)", mat2_sum[63:0]);
        end
        if (mat2_sum[127:64] == 64'h40460A1CAC083127) begin
            $display($time,"ps: Pass! e_12 + f_12 = g_12 (%h)", mat2_sum[127:64]);
        end else begin
            $display($time,"ps: Error! e_12 + f_12 != g_12 (%h)", mat2_sum[127:64]);
        end
        if (mat2_sum[191:128] == 64'h401F000000000000) begin
            $display($time,"ps: Pass! e_13 + f_13 = g_13 (%h)", mat2_sum[191:128]);
        end else begin
            $display($time,"ps: Error! e_13 + f_13 != g_13 (%h)", mat2_sum[191:128]);
        end
        if (mat2_sum[255:192] == 64'h0021FA474C5E1008) begin
            $display($time,"ps: Pass! e_21 + f_21 = g_21 (%h)", mat2_sum[255:192]);
        end else begin
            $display($time,"ps: Error! e_21 + f_21 != g_21 (%h)", mat2_sum[255:192]);
        end
        if (mat2_sum[319:256] == 64'h001D7B6F52D0A0F7) begin
            $display($time,"ps: Pass! e_22 + f_22 = g_22 (%h)", mat2_sum[319:256]);
        end else begin
            $display($time,"ps: Error! e_22 + f_22 != g_22 (%h)", mat2_sum[319:256]);
        end
        if (mat2_sum[383:320] == 64'h404B000000000000) begin
            $display($time,"ps: Pass! e_23 + f_23 = g_23 (%h)", mat2_sum[383:320]);
        end else begin
            $display($time,"ps: Error! e_23 + f_23 != g_23 (%h)", mat2_sum[383:320]);
        end
        if (mat2_sum[447:384] == 64'hC053133333333334) begin
            $display($time,"ps: Pass! e_31 + f_31 = g_31 (%h)", mat2_sum[447:384]);
        end else begin
            $display($time,"ps: Error! e_31 + f_31 != g_31 (%h)", mat2_sum[447:384]);
        end
        if (mat2_sum[511:448] == 64'h000012688B70E62B) begin
            $display($time,"ps: Pass! e_32 + f_32 = g_32 (%h)", mat2_sum[511:448]);
        end else begin
            $display($time,"ps: Error! e_32 + f_32 != g_32 (%h)", mat2_sum[511:448]);
        end
        if (mat2_sum[575:512] == 64'h000003AE8249C7A2) begin
            $display($time,"ps: Pass! e_33 + f_33 = g_33 (%h)", mat2_sum[575:512]);
        end else begin
            $display($time,"ps: Error! e_33 + f_33 != g_33 (%h)", mat2_sum[575:512]);
        end
        #3000000;
        $finish;
    end

    always begin
        #5000;
        clk = ~clk;
    end

endmodule
