`timescale 1ns / 1ns

module rng_uni_tb ();

    reg  clk, rst, mode;
    reg [1023 : 0] init_state;
    wire s_in;
    wire [31 : 0] rng;

    initial begin
        $dumpfile("rng_uni.vcd");
        // $dumpvars(0, rng_uni_tb);
        init_state = 1024'b1001011100111000001000110110101001110000110011111010110101100100001111011110010010110101000000101010100000110101100010101000110011011101110111100101010011000010111010001100000100010011111110100110110000000001001101110010011101111001111111100000000101001101001110000111010111100000100101101010111001110011111100100111010110000100110110010110011101100011011101101001000110111110100111110111100100111101011001001010101111011111111001011100011011000010100100111000010010010000110100111101110011000111101000111110110110001110110110101000000000111101101101001110111100110100111000111000101010110001111010001000001010011010011011010010000101001010011100001010111111111101111100010111000101001100000111011100111100110001110010000001010111111110101010000000100011110011011101111110001100010110111111000010101101011110100111111110001001100111000110111011111000010000000001010101101100011000101011011100100001010010001001111100110101110010000110010111110111010111101001110100100000001110101101011111101001100110111100111100101100000111;
        clk = 1'b0;
        rst = 1'b1;
        mode = 1'b0;
        #30;
        rst = 1'b0;
        mode = 1'b1; // Serial load mode.
        #10240;
        mode = 1'b0; // RNG mode.

        #40000000;
        $finish;
    end

    rng_uni UUT (
    .rng   (rng),
    .s_out (), // Unconnected.
    .s_in  (s_in),
    .ce    (1'b1),
    .mode  (mode),
    .rst   (rst),
    .clk   (clk)
    );

    always @(posedge clk) begin
        if (mode) begin
            init_state <= {init_state[0], init_state[1023 : 1]};
        end else begin
            init_state <= init_state;
            $display("%d", rng);
        end
    end

    assign s_in = init_state[0];

    always begin
        #5 clk = (clk === 1'b0);
    end

endmodule
